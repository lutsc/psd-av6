library ieee;
use ieee.std_logic_1164.all;

entity mdc_top is
end entity;

architecture arch_mdc_top of mdc_top is
begin

end architecture;