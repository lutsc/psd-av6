library ieee;
use ieee.std_logic_1164.all;

entity mdc_datapath is
end entity;

architecture arch_datapath of mdc_datapath is
begin

end architecture;