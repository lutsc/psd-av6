library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity subtractor is port(
  i_CLR_n : in std_logic;
  i_CLK   : in std_logic;
  i_ENA   : in std_logic;
  i_A     : in std_logic_vector(7 downto 0);
  i_B     : in std_logic_vector(7 downto 0);
  o_S     : out std_logic_vector(7 downto 0));
end entity;

architecture arch_subtractor of subtractor is

  signal w_S : std_logic_vector(7 downto 0);

begin
  
  w_S <= std_logic_vector(unsigned(i_A) - unsigned(i_B));

  process(i_CLR_n, i_CLK, i_ENA)
  begin
    if (i_CLR_n = '0') then
      o_S <= (others => '0');
    elsif (rising_edge(i_CLK) and i_ENA = '1') then
      o_S <= w_S;
    end if;
  end process;

end architecture;