library ieee;
use ieee.std_logic_1164.all;

entity mdc_controller is
end entity;

architecture arch_controller of mdc_controller is
begin

end architecture;